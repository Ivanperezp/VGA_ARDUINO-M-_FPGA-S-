module top_vga (
    input  wire        CLOCK_50,  // 50 MHz clock from DE0-CV
    input  wire        RESET_n,   // Active-low reset button
    output wire        VGA_HS,    // Hsync to monitor
    output wire        VGA_VS,    // Vsync to monitor
    output wire [2:0]  VGA_R,     // 3 red bits
    output wire [2:0]  VGA_G,     // 3 green bits
    output wire [1:0]  VGA_B,     // 2 blue bits
    output reg [(ADDR_WIDTH - 1) :0] r_address,
    input [7:0] DATA
);

parameter ADDR_WIDTH = 11;
parameter DIVISION = 16;

//---------------------------------------------------------------------
// 1) Internal signals for PLL and VGA logic
//---------------------------------------------------------------------
wire clk_25MHz;    // 25 MHz clock generated by PLL
wire locked_pll;   // Indicates PLL is stabilized

//---------------------------------------------------------------------
// 2) PLL instance (generated by Quartus IP)
//    File named "prueba_0002.v"
//    Module name "prueba_0002"
//---------------------------------------------------------------------
pll pll_inst (
    .refclk   (CLOCK_50),     // Connect 50 MHz clock
    .rst      (~RESET_n),     // Active-low reset => inverted
    .outclk_0 (clk_25MHz),    // 25 MHz output
    .locked   (locked_pll)
);

//---------------------------------------------------------------------
// 3) Signals for VGA synchronization
//---------------------------------------------------------------------
wire hsync_sig, vsync_sig;
wire video_enable;
wire [9:0] hcount, vcount;

//---------------------------------------------------------------------
// 4) Instantiate VGA synchronization module
//---------------------------------------------------------------------
vga_sync sync_unit (
    .clk_25MHz    (clk_25MHz),
    .reset        (~RESET_n),   // Could use (!locked_pll) for more control -> .reset (~RESET_n | ~locked_pll)
    .hsync        (hsync_sig),
    .vsync        (vsync_sig),
    .video_enable (video_enable),
    .hcount       (hcount),
    .vcount       (vcount)
);

// Connect hsync and vsync signals to top-level outputs
assign VGA_HS = hsync_sig;
assign VGA_VS = vsync_sig;

//---------------------------------------------------------------------
// 5) Color generation logic
//---------------------------------------------------------------------
reg [2:0] color_r;
reg [2:0] color_g;
reg [2:0] color_b;

always @(posedge clk_25MHz) begin
    // While PLL is not locked, we could force black
    if (!locked_pll) begin
        color_r <= 3'b000;
        color_g <= 3'b000;
        color_b <= 3'b000;
    end
    // Outside visible area, paint black
    else if (!video_enable) begin
        color_r <= 3'b000;
        color_g <= 3'b000;
        color_b <= 3'b000;
    end
    // In visible area, generate a simple pattern. Example: half red / half blue
    else begin
        r_address <= (hcount / DIVISION) + (vcount / DIVISION) * (640 / DIVISION);
        
        color_r <= DATA[7:5];
        color_g <= DATA[4:2];
        color_b <= DATA[1:0];
    end
end

// Assign outputs
assign VGA_R = color_r;
assign VGA_G = color_g;
assign VGA_B = color_b;

endmodule